library verilog;
use verilog.vl_types.all;
entity Measure is
end Measure;
